CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
360 300 1 100 10
176 79 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
143654930 0
0
6 Title:
5 Name:
0
0
0
153
13 Logic Switch~
5 995 499 0 10 11
0 136 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -19 8 -11
5 modo1
-15 -26 20 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89649e-315 0
0
13 Logic Switch~
5 154 281 0 10 11
0 142 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
3 set
-8 -26 13 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
41680 0
0
13 Logic Switch~
5 160 498 0 10 11
0 146 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-9 -18 5 -10
4 modo
-12 -26 16 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
41680 2
0
5 4049~
219 181 1188 0 2 22
0 3 4
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U61D
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 61 0
1 U
3421 0 0
2
5.89649e-315 0
0
5 4081~
219 195 1150 0 3 22
0 4 6 5
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U62B
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 62 0
1 U
8157 0 0
2
5.89649e-315 0
0
5 4049~
219 126 1418 0 2 22
0 3 7
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U61C
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 61 0
1 U
5572 0 0
2
41680 3
0
5 4081~
219 139 1381 0 3 22
0 7 9 8
0
0 0 624 90
4 4081
-7 -24 21 -16
4 U62A
17 -5 45 3
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 62 0
1 U
8901 0 0
2
41680 4
0
6 74LS85
106 1062 612 0 14 29
0 11 12 13 14 15 16 17 18 151
152 153 3 10 10
0
0 0 5104 0
5 74F85
-18 -52 17 -44
2 U7
-7 -62 7 -54
0
15 DVCC=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 13 12 10 1 14 11 9 2
3 4 7 6 5 15 13 12 10 1
14 11 9 2 3 4 7 6 5 0
65 0 0 512 1 0 0 0
1 U
7361 0 0
2
41680 5
0
5 4049~
219 302 1518 0 2 22
0 10 3
0
0 0 624 180
4 4049
-7 -24 21 -16
4 U61B
-8 -20 20 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 61 0
1 U
4747 0 0
2
5.89649e-315 5.26354e-315
0
9 CC 7-Seg~
183 473 1634 0 18 19
10 27 28 29 30 31 32 33 34 154
1 1 1 1 1 1 0 1 2
0
0 0 20592 0
5 REDCC
16 -41 51 -33
2 X1
26 -51 40 -43
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.89649e-315 5.30499e-315
0
5 4049~
219 2237 182 0 2 22
0 15 40
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A1F
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 10 0
1 U
3472 0 0
2
5.89649e-315 5.32571e-315
0
5 4049~
219 2335 186 0 2 22
0 18 41
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A1E
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 10 0
1 U
9998 0 0
2
5.89649e-315 5.34643e-315
0
5 4049~
219 2305 185 0 2 22
0 17 44
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A1D
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 10 0
1 U
3536 0 0
2
5.89649e-315 5.3568e-315
0
5 4049~
219 2273 184 0 2 22
0 16 39
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A1C
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 10 0
1 U
4597 0 0
2
5.89649e-315 5.36716e-315
0
8 3-In OR~
219 2819 264 0 4 22
0 78 77 76 27
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U59B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 59 0
1 U
3835 0 0
2
5.89649e-315 5.37752e-315
0
6 74266~
219 2693 311 0 3 22
0 16 18 76
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U60A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 60 0
1 U
3670 0 0
2
5.89649e-315 5.38788e-315
0
5 7415~
219 2703 269 0 4 22
0 40 17 18 77
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U56C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 56 0
1 U
5616 0 0
2
5.89649e-315 5.39306e-315
0
9 2-In AND~
219 2703 226 0 3 22
0 15 44 78
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U58B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 58 0
1 U
9323 0 0
2
5.89649e-315 5.39824e-315
0
8 3-In OR~
219 2822 475 0 4 22
0 70 71 72 28
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U59A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 59 0
1 U
317 0 0
2
5.89649e-315 5.40342e-315
0
9 2-In AND~
219 2432 409 0 3 22
0 44 41 75
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U58A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 58 0
1 U
3108 0 0
2
5.89649e-315 5.4086e-315
0
5 4071~
219 2517 364 0 3 22
0 39 75 70
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U57B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 57 0
1 U
4299 0 0
2
5.89649e-315 5.41378e-315
0
9 2-In AND~
219 2435 461 0 3 22
0 15 44 74
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U54D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 54 0
1 U
9672 0 0
2
5.89649e-315 5.41896e-315
0
9 2-In AND~
219 2435 509 0 3 22
0 15 41 73
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U54C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 54 0
1 U
7876 0 0
2
5.89649e-315 5.42414e-315
0
5 4071~
219 2511 495 0 3 22
0 74 73 71
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U57A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 57 0
1 U
6369 0 0
2
5.89649e-315 5.42933e-315
0
5 7415~
219 2434 558 0 4 22
0 40 17 18 72
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U56B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 56 0
1 U
9172 0 0
2
5.89649e-315 5.43192e-315
0
8 3-In OR~
219 2817 630 0 4 22
0 18 69 68 29
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U52C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 52 0
1 U
7100 0 0
2
5.89649e-315 5.43451e-315
0
6 74266~
219 2554 656 0 3 22
0 16 17 69
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U41D
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 41 0
1 U
3820 0 0
2
5.89649e-315 5.4371e-315
0
6 74266~
219 2555 709 0 3 22
0 15 17 68
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U41C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 41 0
1 U
7678 0 0
2
5.89649e-315 5.43969e-315
0
8 3-In OR~
219 2820 906 0 4 22
0 65 62 59 30
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U52B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 52 0
1 U
961 0 0
2
5.89649e-315 5.44228e-315
0
9 2-In AND~
219 2439 777 0 3 22
0 39 41 66
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U54B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 54 0
1 U
3178 0 0
2
5.89649e-315 5.44487e-315
0
5 7415~
219 2442 825 0 4 22
0 15 16 44 67
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U56A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 56 0
1 U
3409 0 0
2
5.89649e-315 5.44746e-315
0
5 4071~
219 2503 802 0 3 22
0 66 67 65
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U51D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 51 0
1 U
3951 0 0
2
5.89649e-315 5.45005e-315
0
5 7415~
219 2446 882 0 4 22
0 44 16 18 64
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U55C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 55 0
1 U
8885 0 0
2
5.89649e-315 5.45264e-315
0
5 7415~
219 2448 933 0 4 22
0 15 16 18 63
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U55B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 55 0
1 U
3780 0 0
2
5.89649e-315 5.45523e-315
0
5 4071~
219 2516 907 0 3 22
0 64 63 62
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U51C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 51 0
1 U
9265 0 0
2
5.89649e-315 5.45782e-315
0
5 7415~
219 2453 989 0 4 22
0 40 39 17 61
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U55A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 55 0
1 U
9442 0 0
2
5.89649e-315 5.46041e-315
0
5 7415~
219 2455 1049 0 4 22
0 40 17 41 60
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U53C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 53 0
1 U
9424 0 0
2
5.89649e-315 5.463e-315
0
5 4071~
219 2520 1013 0 3 22
0 61 60 59
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U51B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 51 0
1 U
9968 0 0
2
5.89649e-315 5.46559e-315
0
9 2-In AND~
219 2449 1109 0 3 22
0 39 41 58
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U54A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 54 0
1 U
9281 0 0
2
5.89649e-315 5.46818e-315
0
5 7415~
219 2449 1154 0 4 22
0 15 44 41 57
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U53B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 53 0
1 U
8464 0 0
2
5.89649e-315 5.47077e-315
0
5 7415~
219 2448 1201 0 4 22
0 40 17 41 56
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U53A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 53 0
1 U
7168 0 0
2
5.89649e-315 5.47207e-315
0
8 3-In OR~
219 2821 1143 0 4 22
0 58 57 56 31
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U52A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 52 0
1 U
3171 0 0
2
5.89649e-315 5.47336e-315
0
5 7415~
219 2450 1259 0 4 22
0 40 44 41 55
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U50C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 50 0
1 U
4139 0 0
2
5.89649e-315 5.47466e-315
0
5 7415~
219 2452 1308 0 4 22
0 40 16 44 54
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U50B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 50 0
1 U
6435 0 0
2
5.89649e-315 5.47595e-315
0
5 4071~
219 2526 1283 0 3 22
0 55 54 49
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U51A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 51 0
1 U
5283 0 0
2
5.89649e-315 5.47725e-315
0
5 7415~
219 2453 1360 0 4 22
0 15 39 44 53
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U50A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 50 0
1 U
6874 0 0
2
5.89649e-315 5.47854e-315
0
5 7415~
219 2453 1410 0 4 22
0 15 16 17 52
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U35A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 35 0
1 U
5305 0 0
2
5.89649e-315 5.47984e-315
0
5 4071~
219 2529 1384 0 3 22
0 53 52 48
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U34A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 34 0
1 U
34 0 0
2
5.89649e-315 5.48113e-315
0
5 7415~
219 2453 1458 0 4 22
0 16 17 41 51
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U33A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 33 0
1 U
969 0 0
2
5.89649e-315 5.48243e-315
0
5 7415~
219 2454 1504 0 4 22
0 15 17 41 50
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U32A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 32 0
1 U
8402 0 0
2
5.89649e-315 5.48372e-315
0
5 4071~
219 2532 1473 0 3 22
0 51 50 47
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U31A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 31 0
1 U
3751 0 0
2
5.89649e-315 5.48502e-315
0
8 3-In OR~
219 2816 1384 0 4 22
0 49 48 47 32
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U30A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 30 0
1 U
4292 0 0
2
5.89649e-315 5.48631e-315
0
9 2-In AND~
219 2455 1562 0 3 22
0 16 44 46
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U29A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
6118 0 0
2
5.89649e-315 5.48761e-315
0
9 2-In AND~
219 2457 1608 0 3 22
0 15 44 45
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U27A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 27 0
1 U
34 0 0
2
5.89649e-315 5.4889e-315
0
5 4071~
219 2526 1582 0 3 22
0 46 45 38
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U26A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 26 0
1 U
6357 0 0
2
5.89649e-315 5.4902e-315
0
9 2-In AND~
219 2457 1654 0 3 22
0 15 16 43
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 48 0
1 U
319 0 0
2
5.89649e-315 5.49149e-315
0
5 4071~
219 2521 1678 0 3 22
0 43 42 37
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U25A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 25 0
1 U
3976 0 0
2
5.89649e-315 5.49279e-315
0
5 7415~
219 2459 1704 0 4 22
0 16 17 41 42
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U24A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 24 0
1 U
7634 0 0
2
5.89649e-315 5.49408e-315
0
5 7415~
219 2459 1754 0 4 22
0 40 39 17 36
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U49C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 49 0
1 U
523 0 0
2
5.89649e-315 5.49538e-315
0
8 3-In OR~
219 2826 1632 0 4 22
0 38 37 36 33
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U23A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 23 0
1 U
6748 0 0
2
5.89649e-315 5.49667e-315
0
9 2-In AND~
219 2540 1813 0 3 22
0 15 35 34
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 48 0
1 U
6901 0 0
2
5.89649e-315 5.49797e-315
0
5 4071~
219 2443 1837 0 3 22
0 16 17 35
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U47D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 47 0
1 U
842 0 0
2
5.89649e-315 5.49926e-315
0
5 4071~
219 1402 1836 0 3 22
0 12 13 79
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U47C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 47 0
1 U
3277 0 0
2
5.89649e-315 5.50056e-315
0
9 2-In AND~
219 1499 1812 0 3 22
0 11 79 26
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 48 0
1 U
4212 0 0
2
5.89649e-315 5.50185e-315
0
8 3-In OR~
219 1785 1631 0 4 22
0 82 81 80 25
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U40C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 40 0
1 U
4720 0 0
2
5.89649e-315 5.50315e-315
0
5 7415~
219 1418 1753 0 4 22
0 84 83 13 80
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U49B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 49 0
1 U
5551 0 0
2
5.89649e-315 5.50444e-315
0
5 7415~
219 1418 1703 0 4 22
0 12 13 85 86
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U49A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 49 0
1 U
6986 0 0
2
5.89649e-315 5.50574e-315
0
5 4071~
219 1480 1677 0 3 22
0 87 86 81
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U47B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 47 0
1 U
8745 0 0
2
5.89649e-315 5.50703e-315
0
9 2-In AND~
219 1416 1653 0 3 22
0 11 12 87
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U48A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 48 0
1 U
9592 0 0
2
5.89649e-315 5.50833e-315
0
5 4071~
219 1485 1581 0 3 22
0 90 89 82
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U47A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 47 0
1 U
8748 0 0
2
5.89649e-315 5.50963e-315
0
9 2-In AND~
219 1416 1607 0 3 22
0 11 88 89
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U42D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 42 0
1 U
7168 0 0
2
5.89649e-315 5.51092e-315
0
9 2-In AND~
219 1414 1561 0 3 22
0 12 88 90
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U42C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 42 0
1 U
631 0 0
2
5.89649e-315 5.51222e-315
0
8 3-In OR~
219 1775 1383 0 4 22
0 93 92 91 24
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U40B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 40 0
1 U
9466 0 0
2
5.89649e-315 5.51286e-315
0
5 4071~
219 1491 1472 0 3 22
0 95 94 91
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U44D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 44 0
1 U
3266 0 0
2
5.89649e-315 5.51351e-315
0
5 7415~
219 1413 1503 0 4 22
0 11 13 85 94
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U46C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 46 0
1 U
7693 0 0
2
5.89649e-315 5.51416e-315
0
5 7415~
219 1412 1457 0 4 22
0 12 13 85 95
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U46B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 46 0
1 U
3723 0 0
2
5.89649e-315 5.51481e-315
0
5 4071~
219 1488 1383 0 3 22
0 97 96 92
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U44C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 44 0
1 U
3440 0 0
2
5.89649e-315 5.51545e-315
0
5 7415~
219 1412 1409 0 4 22
0 11 12 13 96
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U46A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 46 0
1 U
6263 0 0
2
5.89649e-315 5.5161e-315
0
5 7415~
219 1412 1359 0 4 22
0 11 83 88 97
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U45C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 45 0
1 U
4900 0 0
2
5.89649e-315 5.51675e-315
0
5 4071~
219 1485 1282 0 3 22
0 99 98 93
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U44B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 44 0
1 U
8783 0 0
2
5.89649e-315 5.5174e-315
0
5 7415~
219 1411 1307 0 4 22
0 84 12 88 98
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U45B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 45 0
1 U
3221 0 0
2
5.89649e-315 5.51804e-315
0
5 7415~
219 1409 1258 0 4 22
0 84 88 85 99
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U45A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 45 0
1 U
3215 0 0
2
5.89649e-315 5.51869e-315
0
8 3-In OR~
219 1780 1142 0 4 22
0 102 101 100 23
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U40A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 40 0
1 U
7903 0 0
2
5.89649e-315 5.51934e-315
0
5 7415~
219 1407 1200 0 4 22
0 84 13 85 100
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U22A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 22 0
1 U
7121 0 0
2
5.89649e-315 5.51999e-315
0
5 7415~
219 1408 1153 0 4 22
0 11 88 85 101
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U21A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 21 0
1 U
4484 0 0
2
5.89649e-315 5.52063e-315
0
9 2-In AND~
219 1408 1108 0 3 22
0 83 85 102
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U42B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 42 0
1 U
5996 0 0
2
5.89649e-315 5.52128e-315
0
5 4071~
219 1479 1012 0 3 22
0 105 104 103
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U44A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 44 0
1 U
7804 0 0
2
5.89649e-315 5.52193e-315
0
5 7415~
219 1414 1048 0 4 22
0 84 13 85 104
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U19A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 19 0
1 U
5523 0 0
2
5.89649e-315 5.52258e-315
0
5 7415~
219 1412 988 0 4 22
0 84 83 13 105
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 18 0
1 U
3330 0 0
2
5.89649e-315 5.52322e-315
0
5 4071~
219 1475 906 0 3 22
0 108 107 106
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U15D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 15 0
1 U
3465 0 0
2
5.89649e-315 5.52387e-315
0
5 7415~
219 1407 932 0 4 22
0 11 12 14 107
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 43 0
1 U
8396 0 0
2
5.89649e-315 5.52452e-315
0
5 7415~
219 1405 881 0 4 22
0 88 12 14 108
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 43 0
1 U
3685 0 0
2
5.89649e-315 5.52517e-315
0
5 4071~
219 1462 801 0 3 22
0 110 111 109
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U15C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 15 0
1 U
7849 0 0
2
5.89649e-315 5.52581e-315
0
5 7415~
219 1401 824 0 4 22
0 11 12 88 111
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U43A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 43 0
1 U
6343 0 0
2
5.89649e-315 5.52646e-315
0
9 2-In AND~
219 1398 776 0 3 22
0 83 85 110
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U42A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 42 0
1 U
7376 0 0
2
5.89649e-315 5.52711e-315
0
8 3-In OR~
219 1779 905 0 4 22
0 109 106 103 22
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U17A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 17 0
1 U
9156 0 0
2
5.89649e-315 5.52776e-315
0
6 74266~
219 1514 708 0 3 22
0 11 13 112
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U41B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 41 0
1 U
5776 0 0
2
5.89649e-315 5.52841e-315
0
6 74266~
219 1513 655 0 3 22
0 12 13 113
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U41A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
7207 0 0
2
5.89649e-315 5.52905e-315
0
8 3-In OR~
219 1776 629 0 4 22
0 14 113 112 21
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U20A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 20 0
1 U
4459 0 0
2
5.89649e-315 5.5297e-315
0
5 7415~
219 1393 557 0 4 22
0 84 13 14 116
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U16A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 16 0
1 U
3760 0 0
2
5.89649e-315 5.53035e-315
0
5 4071~
219 1470 494 0 3 22
0 118 117 115
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U15B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 15 0
1 U
754 0 0
2
5.89649e-315 5.531e-315
0
9 2-In AND~
219 1394 508 0 3 22
0 11 85 117
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U39D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 39 0
1 U
9767 0 0
2
5.89649e-315 5.53164e-315
0
9 2-In AND~
219 1394 460 0 3 22
0 11 88 118
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U39C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 39 0
1 U
7978 0 0
2
5.89649e-315 5.53229e-315
0
5 4071~
219 1476 363 0 3 22
0 83 119 114
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U15A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 15 0
1 U
3142 0 0
2
5.89649e-315 5.53294e-315
0
9 2-In AND~
219 1391 408 0 3 22
0 88 85 119
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U39B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 39 0
1 U
3284 0 0
2
5.89649e-315 5.53359e-315
0
8 3-In OR~
219 1781 474 0 4 22
0 114 115 116 20
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U36C
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 36 0
1 U
659 0 0
2
5.89649e-315 5.53423e-315
0
5 4030~
219 600 797 0 3 22
0 145 144 120
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U38A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 38 0
1 U
3800 0 0
2
41680 6
0
5 7422~
219 218 1441 0 5 22
0 121 124 123 122 9
0
0 0 624 512
6 74LS22
-21 -28 21 -20
4 U37A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 37 0
1 U
6792 0 0
2
41680 7
0
14 Logic Display~
6 68 1083 0 1 2
13 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 OVERF
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3701 0 0
2
41680 8
0
14 Logic Display~
6 131 1043 0 1 2
22 8
0
0 0 53872 0
6 100MEG
2 -16 44 -8
6 PERDEU
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6316 0 0
2
41680 9
0
14 Logic Display~
6 193 1004 0 1 2
12 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
6 GANHOU
-21 -21 21 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8734 0 0
2
41680 10
0
9 4-In AND~
219 304 1339 0 5 22
0 121 123 124 122 6
0
0 0 624 512
6 74LS21
-21 -28 21 -20
4 U11A
-16 -28 12 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 12 0
1 U
7988 0 0
2
41680 11
0
6 74266~
219 465 1209 0 3 22
0 132 128 121
0
0 0 624 512
7 74LS266
-24 -24 25 -16
4 U28C
1 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
3217 0 0
2
41680 12
0
6 74266~
219 466 1298 0 3 22
0 131 127 123
0
0 0 624 512
7 74LS266
-24 -24 25 -16
4 U28D
1 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
3965 0 0
2
41680 13
0
6 74266~
219 468 1386 0 3 22
0 130 126 124
0
0 0 624 512
7 74LS266
-24 -24 25 -16
3 U9A
4 -25 25 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8239 0 0
2
41680 14
0
6 74266~
219 469 1461 0 3 22
0 129 125 122
0
0 0 624 512
7 74LS266
-24 -24 25 -16
4 U10A
1 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
828 0 0
2
41680 15
0
8 Hex Key~
166 678 1083 0 11 12
0 129 130 131 132 0 0 0 0 0
5 53
0
0 0 4656 0
0
7 Entrada
-25 -34 24 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
6187 0 0
2
41680 16
0
9 2-In AND~
219 1662 225 0 3 22
0 11 88 135
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7107 0 0
2
5.89649e-315 5.53488e-315
0
5 7415~
219 1662 268 0 4 22
0 84 13 14 134
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 U12A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 11 0
1 U
6433 0 0
2
5.89649e-315 5.53553e-315
0
6 74266~
219 1652 310 0 3 22
0 12 14 133
0
0 0 624 0
7 74LS266
-24 -24 25 -16
4 U13A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
8559 0 0
2
5.89649e-315 5.53618e-315
0
8 3-In OR~
219 1778 263 0 4 22
0 135 134 133 19
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 14 0
1 U
3674 0 0
2
5.89649e-315 5.53682e-315
0
5 4049~
219 1231 127 0 2 22
0 12 83
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A13
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 9 0
1 U
5697 0 0
2
5.89649e-315 5.53747e-315
0
5 4049~
219 1262 129 0 2 22
0 13 88
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A14
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 10 0
1 U
3805 0 0
2
5.89649e-315 5.53812e-315
0
5 4049~
219 1294 129 0 2 22
0 14 85
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A15
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 10 0
1 U
5219 0 0
2
5.89649e-315 5.53877e-315
0
5 4049~
219 1197 127 0 2 22
0 11 84
0
0 0 112 270
4 4049
-7 -24 21 -16
3 A16
-4 -34 17 -26
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 9 0
1 U
3795 0 0
2
5.89649e-315 5.53941e-315
0
9 CC 7-Seg~
183 225 1633 0 18 19
10 19 20 21 22 23 24 25 26 155
1 1 1 0 0 1 1 0 2
0
0 0 20592 0
5 REDCC
16 -41 51 -33
2 X2
26 -51 40 -43
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3637 0 0
2
5.89649e-315 5.54006e-315
0
5 4049~
219 922 528 0 2 22
0 18 137
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 9 0
1 U
3226 0 0
2
5.89649e-315 5.54071e-315
0
5 4049~
219 921 457 0 2 22
0 16 139
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 9 0
1 U
6966 0 0
2
5.89649e-315 5.54136e-315
0
5 4049~
219 921 490 0 2 22
0 17 138
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
9796 0 0
2
5.89649e-315 5.542e-315
0
5 4049~
219 921 423 0 2 22
0 15 140
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
5952 0 0
2
5.89649e-315 5.54265e-315
0
6 74LS83
105 1048 448 0 14 29
0 11 12 13 14 140 139 138 137 136
128 127 126 125 156
0
0 0 4848 0
5 74F83
-18 -60 17 -52
3 ULA
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3649 0 0
2
5.89649e-315 5.5433e-315
0
14 Logic Display~
6 687 579 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3716 0 0
2
41680 17
0
14 Logic Display~
6 730 578 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4797 0 0
2
41680 18
0
14 Logic Display~
6 775 579 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4681 0 0
2
41680 19
0
14 Logic Display~
6 803 579 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9730 0 0
2
41680 20
0
2 +V
167 252 755 0 1 3
0 141
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9874 0 0
2
41680 21
0
6 JK RN~
219 816 800 0 6 22
0 17 2 17 141 157 18
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
364 0 0
2
41680 22
0
6 JK RN~
219 706 801 0 6 22
0 143 2 120 141 158 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
3656 0 0
2
41680 23
0
6 JK RN~
219 493 787 0 6 22
0 15 2 15 141 145 16
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 1 0
1 U
3131 0 0
2
41680 24
0
6 JK RN~
219 381 778 0 6 22
0 141 2 141 141 144 15
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 1 0
1 U
6772 0 0
2
41680 25
0
14 Logic Display~
6 790 88 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9557 0 0
2
41680 26
0
14 Logic Display~
6 835 94 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5789 0 0
2
41680 27
0
14 Logic Display~
6 883 95 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7328 0 0
2
41680 28
0
14 Logic Display~
6 935 95 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4799 0 0
2
41680 29
0
9 2-In AND~
219 311 427 0 3 22
0 147 146 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
9196 0 0
2
41680 33
0
7 Pulser~
4 130 399 0 10 12
0 159 160 147 161 0 0 16 16 1
7
0
0 0 4656 0
0
5 Pulso
-17 -28 18 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3857 0 0
2
41680 34
0
6 74112~
219 253 270 0 7 32
0 142 148 2 148 141 162 11
0
0 0 4720 180
7 74LS112
-3 -60 46 -52
3 U2B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 2 0
1 U
7125 0 0
2
41680 35
0
6 74112~
219 441 270 0 7 32
0 142 149 2 149 141 163 12
0
0 0 4720 180
7 74LS112
-3 -60 46 -52
3 U2A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 1 2 0
1 U
3641 0 0
2
41680 36
0
6 74112~
219 617 270 0 7 32
0 142 14 2 14 141 164 13
0
0 0 4720 180
7 74LS112
-3 -60 46 -52
3 U1B
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0
65 0 0 512 2 2 1 0
1 U
9821 0 0
2
41680 37
0
2 +V
167 925 226 0 1 3
0 150
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3187 0 0
2
41680 38
0
5 4073~
219 325 104 0 4 22
0 12 13 14 148
0
0 0 624 180
4 4073
-7 -24 21 -16
3 U4A
-13 -25 8 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
762 0 0
2
41680 39
0
9 2-In AND~
219 595 144 0 3 22
0 13 14 149
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U3A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
39 0 0
2
41680 40
0
6 74112~
219 788 271 0 7 32
0 142 150 2 150 141 165 14
0
0 0 4720 180
7 74LS112
-3 -60 46 -52
3 U1A
21 -63 42 -55
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
22

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 1872418908
65 0 0 512 2 1 1 0
1 U
9450 0 0
2
41680 41
0
375
3 0 2 0 0 8192 0 145 0 0 360 3
332 427
332 425
426 425
1 0 3 0 0 4096 0 4 0 0 20 2
184 1206
68 1206
2 1 4 0 0 4224 0 4 5 0 0 3
184 1170
184 1171
185 1171
3 1 5 0 0 12416 0 5 111 0 0 4
194 1126
194 1127
193 1127
193 1022
5 2 6 0 0 8320 0 112 5 0 0 3
279 1339
203 1339
203 1171
1 0 3 0 0 0 0 6 0 0 20 2
129 1436
68 1436
2 1 7 0 0 4224 0 6 7 0 0 2
129 1400
129 1402
3 1 8 0 0 4224 0 7 110 0 0 4
138 1357
138 1080
131 1080
131 1061
2 5 9 0 0 8320 0 7 108 0 0 3
147 1402
147 1441
193 1441
2 0 3 0 0 8192 0 9 0 0 20 4
287 1518
83 1518
83 1105
68 1105
14 0 10 0 0 8192 0 8 0 0 21 3
1094 648
1094 653
1168 653
0 1 11 0 0 4096 0 0 8 321 0 3
1009 400
1009 585
1030 585
0 2 12 0 0 4096 0 0 8 320 0 3
996 419
996 594
1030 594
0 3 13 0 0 4096 0 0 8 319 0 3
991 430
991 603
1030 603
0 4 14 0 0 4096 0 0 8 318 0 3
977 439
977 612
1030 612
0 5 15 0 0 12288 0 0 8 158 0 4
950 632
982 632
982 621
1030 621
0 6 16 0 0 12288 0 0 8 156 0 4
958 646
989 646
989 630
1030 630
0 7 17 0 0 4096 0 0 8 153 0 4
965 669
1010 669
1010 639
1030 639
0 8 18 0 0 4096 0 0 8 155 0 3
972 694
1030 694
1030 648
12 1 3 0 0 16512 0 8 109 0 0 6
1094 630
1094 628
1173 628
1173 1538
68 1538
68 1101
13 1 10 0 0 12416 0 8 9 0 0 5
1094 639
1094 641
1168 641
1168 1518
323 1518
4 1 19 0 0 20608 0 121 126 0 0 7
1811 263
1961 263
1961 16
3025 16
3025 2071
204 2071
204 1669
4 2 20 0 0 20608 0 106 126 0 0 7
1814 474
1970 474
1970 23
3017 23
3017 2058
210 2058
210 1669
4 3 21 0 0 20608 0 99 126 0 0 7
1809 629
1978 629
1978 31
3005 31
3005 2046
216 2046
216 1669
4 4 22 0 0 20608 0 96 126 0 0 7
1812 905
1990 905
1990 41
2995 41
2995 2037
222 2037
222 1669
4 5 23 0 0 20608 0 83 126 0 0 7
1813 1142
1998 1142
1998 50
2987 50
2987 2026
228 2026
228 1669
4 6 24 0 0 20608 0 73 126 0 0 7
1808 1383
2007 1383
2007 61
2978 61
2978 2017
234 2017
234 1669
4 7 25 0 0 20608 0 65 126 0 0 7
1818 1631
2014 1631
2014 68
2970 68
2970 2009
240 2009
240 1669
3 8 26 0 0 20608 0 64 126 0 0 7
1520 1812
2022 1812
2022 77
2962 77
2962 2002
246 2002
246 1669
1 0 18 0 0 4096 0 12 0 0 155 2
2338 168
2338 95
1 0 17 0 0 4096 0 13 0 0 153 2
2308 167
2308 105
1 0 16 0 0 4096 0 14 0 0 156 2
2276 166
2276 114
1 0 15 0 0 0 0 11 0 0 158 2
2240 164
2240 125
4 1 27 0 0 12416 0 15 10 0 0 5
2852 264
2926 264
2926 1965
452 1965
452 1670
4 2 28 0 0 12416 0 19 10 0 0 5
2855 475
2920 475
2920 1955
458 1955
458 1670
4 3 29 0 0 12416 0 26 10 0 0 5
2850 630
2909 630
2909 1944
464 1944
464 1670
4 4 30 0 0 12416 0 29 10 0 0 5
2853 906
2899 906
2899 1935
470 1935
470 1670
4 5 31 0 0 12416 0 42 10 0 0 5
2854 1143
2890 1143
2890 1927
476 1927
476 1670
4 6 32 0 0 12416 0 52 10 0 0 5
2849 1384
2883 1384
2883 1922
482 1922
482 1670
4 7 33 0 0 12416 0 60 10 0 0 5
2859 1632
2875 1632
2875 1912
488 1912
488 1670
3 8 34 0 0 12416 0 61 10 0 0 5
2561 1813
2572 1813
2572 1903
494 1903
494 1670
0 1 15 0 0 8192 0 0 61 56 0 3
2258 1644
2258 1804
2516 1804
3 2 35 0 0 8320 0 62 61 0 0 3
2476 1837
2476 1822
2516 1822
0 2 17 0 0 8192 0 0 62 49 0 3
2323 1763
2323 1846
2430 1846
0 1 16 0 0 8192 0 0 62 54 0 3
2295 1694
2295 1828
2430 1828
3 4 36 0 0 12416 0 60 59 0 0 4
2813 1641
2768 1641
2768 1754
2480 1754
3 2 37 0 0 4224 0 57 60 0 0 4
2554 1678
2752 1678
2752 1632
2814 1632
3 1 38 0 0 4224 0 55 60 0 0 4
2559 1582
2805 1582
2805 1623
2813 1623
0 3 17 0 0 8192 0 0 59 53 0 3
2323 1702
2323 1763
2435 1763
0 2 39 0 0 4096 0 0 59 80 0 3
2275 1358
2275 1754
2435 1754
0 1 40 0 0 4224 0 0 59 90 0 3
2241 1298
2241 1745
2435 1745
0 3 41 0 0 4096 0 0 58 69 0 3
2338 1513
2338 1713
2435 1713
0 2 17 0 0 4096 0 0 58 71 0 3
2323 1502
2323 1704
2435 1704
0 1 16 0 0 8192 0 0 58 55 0 3
2295 1663
2295 1695
2435 1695
0 2 16 0 0 0 0 0 56 62 0 3
2295 1556
2295 1663
2433 1663
0 1 15 0 0 0 0 0 56 60 0 3
2258 1598
2258 1645
2433 1645
4 2 42 0 0 4224 0 58 57 0 0 3
2480 1704
2508 1704
2508 1687
3 1 43 0 0 4224 0 56 57 0 0 3
2478 1654
2508 1654
2508 1669
0 2 44 0 0 8192 0 0 54 61 0 3
2309 1571
2309 1617
2433 1617
0 1 15 0 0 0 0 0 54 73 0 3
2258 1494
2258 1599
2433 1599
0 2 44 0 0 4096 0 0 53 78 0 3
2309 1369
2309 1571
2431 1571
0 1 16 0 0 0 0 0 53 74 0 4
2295 1449
2295 1556
2431 1556
2431 1553
3 2 45 0 0 4224 0 54 55 0 0 4
2478 1608
2509 1608
2509 1591
2513 1591
3 1 46 0 0 4224 0 53 55 0 0 4
2476 1562
2509 1562
2509 1573
2513 1573
3 0 41 0 0 0 0 43 0 0 70 2
2426 1268
2338 1268
3 3 47 0 0 4224 0 51 52 0 0 4
2565 1473
2782 1473
2782 1393
2803 1393
3 2 48 0 0 4224 0 48 52 0 0 2
2562 1384
2804 1384
3 1 49 0 0 4224 0 45 52 0 0 4
2559 1283
2781 1283
2781 1375
2803 1375
0 3 41 0 0 0 0 0 50 70 0 3
2338 1465
2338 1513
2430 1513
0 3 41 0 0 4096 0 0 49 97 0 3
2338 1209
2338 1467
2429 1467
0 2 17 0 0 0 0 0 50 72 0 3
2323 1458
2323 1504
2430 1504
0 2 17 0 0 0 0 0 49 77 0 3
2323 1419
2323 1458
2429 1458
0 1 15 0 0 0 0 0 50 81 0 3
2258 1400
2258 1495
2430 1495
0 1 16 0 0 0 0 0 49 79 0 3
2295 1410
2295 1449
2429 1449
2 4 50 0 0 12416 0 51 50 0 0 4
2519 1482
2511 1482
2511 1504
2475 1504
4 1 51 0 0 4224 0 49 51 0 0 4
2474 1458
2510 1458
2510 1464
2519 1464
0 3 17 0 0 4096 0 0 47 95 0 3
2323 1201
2323 1419
2429 1419
0 3 44 0 0 0 0 0 46 88 0 3
2309 1317
2309 1369
2429 1369
0 2 16 0 0 0 0 0 47 87 0 3
2295 1308
2295 1410
2429 1410
0 2 39 0 0 0 0 0 46 102 0 3
2275 1098
2275 1360
2429 1360
0 1 15 0 0 0 0 0 47 82 0 3
2258 1347
2258 1401
2429 1401
0 1 15 0 0 0 0 0 46 100 0 3
2258 1143
2258 1351
2429 1351
4 2 52 0 0 4224 0 47 48 0 0 4
2474 1410
2507 1410
2507 1393
2516 1393
4 1 53 0 0 4224 0 46 48 0 0 4
2474 1360
2506 1360
2506 1375
2516 1375
4 2 54 0 0 4224 0 44 45 0 0 4
2473 1308
2498 1308
2498 1292
2513 1292
4 1 55 0 0 4224 0 43 45 0 0 4
2471 1259
2500 1259
2500 1274
2513 1274
0 2 16 0 0 4096 0 0 44 117 0 3
2295 933
2295 1308
2428 1308
0 3 44 0 0 0 0 0 44 89 0 3
2309 1257
2309 1317
2428 1317
0 2 44 0 0 0 0 0 43 99 0 3
2309 1157
2309 1259
2426 1259
0 1 40 0 0 0 0 0 44 91 0 3
2241 1250
2241 1299
2428 1299
0 1 40 0 0 0 0 0 43 96 0 3
2241 1190
2241 1250
2426 1250
4 3 56 0 0 4224 0 41 42 0 0 4
2469 1201
2799 1201
2799 1152
2808 1152
4 2 57 0 0 4224 0 40 42 0 0 4
2470 1154
2662 1154
2662 1143
2809 1143
3 1 58 0 0 4224 0 39 42 0 0 4
2470 1109
2798 1109
2798 1134
2808 1134
0 2 17 0 0 0 0 0 41 106 0 3
2323 1049
2323 1201
2424 1201
0 1 40 0 0 0 0 0 41 107 0 3
2241 1040
2241 1192
2424 1192
0 3 41 0 0 0 0 0 41 98 0 3
2338 1163
2338 1210
2424 1210
0 3 41 0 0 0 0 0 40 101 0 3
2338 1118
2338 1163
2425 1163
0 2 44 0 0 4096 0 0 40 119 0 4
2309 871
2309 1157
2425 1157
2425 1154
0 1 15 0 0 0 0 0 40 118 0 3
2258 922
2258 1145
2425 1145
0 2 41 0 0 0 0 0 39 105 0 3
2338 1058
2338 1118
2425 1118
0 1 39 0 0 0 0 0 39 109 0 3
2275 989
2275 1100
2425 1100
0 3 18 0 0 0 0 0 34 104 0 3
2357 891
2357 942
2424 942
0 3 18 0 0 4096 0 0 33 135 0 3
2357 620
2357 891
2422 891
0 3 41 0 0 4224 0 0 37 127 0 3
2338 786
2338 1058
2431 1058
0 2 17 0 0 0 0 0 37 108 0 3
2323 998
2323 1049
2431 1049
0 1 40 0 0 0 0 0 37 110 0 3
2241 980
2241 1040
2431 1040
0 3 17 0 0 4096 0 0 36 132 0 3
2323 718
2323 998
2429 998
0 2 39 0 0 0 0 0 36 128 0 3
2275 767
2275 989
2429 989
0 1 40 0 0 0 0 0 36 141 0 3
2241 548
2241 980
2429 980
3 3 59 0 0 4224 0 38 29 0 0 4
2553 1013
2792 1013
2792 915
2807 915
4 2 60 0 0 4224 0 37 38 0 0 3
2476 1049
2507 1049
2507 1022
4 1 61 0 0 4224 0 36 38 0 0 3
2474 989
2507 989
2507 1004
3 2 62 0 0 4224 0 35 29 0 0 3
2549 907
2808 907
2808 906
4 2 63 0 0 4224 0 34 35 0 0 3
2469 933
2503 933
2503 916
4 1 64 0 0 4224 0 33 35 0 0 3
2467 882
2503 882
2503 898
0 2 16 0 0 0 0 0 34 120 0 3
2295 882
2295 933
2424 933
0 1 15 0 0 0 0 0 34 126 0 3
2258 815
2258 924
2424 924
0 1 44 0 0 0 0 0 33 124 0 3
2309 833
2309 873
2422 873
0 2 16 0 0 0 0 0 33 125 0 3
2295 825
2295 882
2422 882
3 1 65 0 0 4224 0 32 29 0 0 4
2536 802
2791 802
2791 897
2807 897
3 1 66 0 0 4224 0 30 32 0 0 4
2460 777
2483 777
2483 793
2490 793
4 2 67 0 0 4224 0 31 32 0 0 4
2463 825
2484 825
2484 811
2490 811
0 3 44 0 0 4096 0 0 31 145 0 3
2309 470
2309 834
2418 834
0 2 16 0 0 0 0 0 31 134 0 3
2295 647
2295 825
2418 825
0 1 15 0 0 0 0 0 31 131 0 3
2258 703
2258 816
2418 816
0 2 41 0 0 0 0 0 30 144 0 3
2338 518
2338 786
2415 786
0 1 39 0 0 4224 0 0 30 150 0 3
2275 355
2275 768
2415 768
3 3 68 0 0 12416 0 26 28 0 0 4
2804 639
2764 639
2764 709
2594 709
3 2 69 0 0 4224 0 27 26 0 0 4
2593 656
2756 656
2756 630
2805 630
0 1 15 0 0 8192 0 0 28 146 0 4
2258 498
2258 703
2539 703
2539 700
2 0 17 0 0 0 0 28 0 0 133 3
2539 718
2323 718
2323 665
0 2 17 0 0 0 0 0 27 140 0 3
2323 558
2323 665
2538 665
0 1 16 0 0 0 0 0 27 156 0 3
2292 302
2292 647
2538 647
0 1 18 0 0 8192 0 0 26 139 0 3
2357 620
2357 621
2804 621
3 1 70 0 0 4224 0 21 19 0 0 4
2550 364
2775 364
2775 466
2809 466
3 2 71 0 0 4224 0 24 19 0 0 4
2544 495
2774 495
2774 475
2810 475
4 3 72 0 0 4224 0 25 19 0 0 4
2455 558
2804 558
2804 484
2809 484
0 3 18 0 0 0 0 0 25 155 0 5
2357 320
2357 620
2357 620
2357 567
2410 567
0 2 17 0 0 4096 0 0 25 153 0 3
2323 268
2323 558
2410 558
0 1 40 0 0 0 0 0 25 154 0 3
2241 260
2241 549
2410 549
3 2 73 0 0 4224 0 23 24 0 0 4
2456 509
2494 509
2494 504
2498 504
3 1 74 0 0 4224 0 22 24 0 0 3
2456 461
2498 461
2498 486
0 2 41 0 0 0 0 0 23 148 0 3
2338 463
2338 518
2411 518
0 2 44 0 0 0 0 0 22 149 0 3
2306 445
2306 470
2411 470
0 1 15 0 0 0 0 0 23 147 0 3
2258 498
2258 500
2411 500
0 1 15 0 0 0 0 0 22 158 0 5
2258 217
2258 498
2258 498
2258 452
2411 452
2 2 41 0 0 0 0 12 20 0 0 5
2338 204
2338 463
2338 463
2338 418
2408 418
0 1 44 0 0 0 0 0 20 157 0 5
2306 235
2306 445
2306 445
2306 400
2408 400
1 2 39 0 0 0 0 21 14 0 0 5
2504 355
2275 355
2275 355
2276 355
2276 202
3 2 75 0 0 8320 0 20 21 0 0 3
2453 409
2453 373
2504 373
0 3 18 0 0 0 0 0 17 155 0 3
2357 281
2679 281
2679 278
0 2 17 0 0 16512 0 0 17 313 0 8
880 588
965 588
965 1871
2072 1871
2072 105
2323 105
2323 269
2679 269
2 1 40 0 0 0 0 11 17 0 0 3
2240 200
2240 260
2679 260
0 2 18 0 0 16512 0 0 16 294 0 8
900 574
972 574
972 1864
2061 1864
2061 95
2357 95
2357 320
2677 320
0 1 16 0 0 16512 0 0 16 312 0 8
870 604
958 604
958 1880
2080 1880
2080 114
2292 114
2292 302
2677 302
2 2 44 0 0 16512 0 13 18 0 0 5
2308 203
2308 235
2306 235
2306 235
2679 235
0 1 15 0 0 16512 0 0 18 311 0 8
860 619
950 619
950 1889
2088 1889
2088 125
2258 125
2258 217
2679 217
3 3 76 0 0 4224 0 16 15 0 0 3
2732 311
2806 311
2806 273
4 2 77 0 0 4224 0 17 15 0 0 3
2724 269
2807 269
2807 264
3 1 78 0 0 4224 0 18 15 0 0 3
2724 226
2806 226
2806 255
0 1 11 0 0 8192 0 0 64 176 0 3
1217 1643
1217 1803
1475 1803
3 2 79 0 0 8320 0 63 64 0 0 3
1435 1836
1435 1821
1475 1821
0 2 13 0 0 0 0 0 63 169 0 3
1282 1762
1282 1845
1389 1845
0 1 12 0 0 0 0 0 63 174 0 3
1254 1693
1254 1827
1389 1827
3 4 80 0 0 12416 0 65 66 0 0 4
1772 1640
1727 1640
1727 1753
1439 1753
3 2 81 0 0 4224 0 68 65 0 0 4
1513 1677
1711 1677
1711 1631
1773 1631
3 1 82 0 0 4224 0 70 65 0 0 4
1518 1581
1764 1581
1764 1622
1772 1622
0 3 13 0 0 0 0 0 66 173 0 3
1282 1701
1282 1762
1394 1762
0 2 83 0 0 4096 0 0 66 200 0 3
1234 1357
1234 1753
1394 1753
0 1 84 0 0 4224 0 0 66 210 0 3
1200 1297
1200 1744
1394 1744
0 3 85 0 0 4096 0 0 67 189 0 3
1297 1512
1297 1712
1394 1712
0 2 13 0 0 4096 0 0 67 191 0 3
1282 1501
1282 1703
1394 1703
0 1 12 0 0 0 0 0 67 175 0 3
1254 1662
1254 1694
1394 1694
0 2 12 0 0 0 0 0 69 182 0 3
1254 1555
1254 1662
1392 1662
0 1 11 0 0 0 0 0 69 180 0 3
1217 1597
1217 1644
1392 1644
4 2 86 0 0 4224 0 67 68 0 0 3
1439 1703
1467 1703
1467 1686
3 1 87 0 0 4224 0 69 68 0 0 3
1437 1653
1467 1653
1467 1668
0 2 88 0 0 8192 0 0 71 181 0 3
1268 1570
1268 1616
1392 1616
0 1 11 0 0 0 0 0 71 193 0 3
1217 1493
1217 1598
1392 1598
0 2 88 0 0 4096 0 0 72 198 0 3
1268 1368
1268 1570
1390 1570
0 1 12 0 0 0 0 0 72 194 0 4
1254 1448
1254 1555
1390 1555
1390 1552
3 2 89 0 0 4224 0 71 70 0 0 4
1437 1607
1468 1607
1468 1590
1472 1590
3 1 90 0 0 4224 0 72 70 0 0 4
1435 1561
1468 1561
1468 1572
1472 1572
3 0 85 0 0 0 0 82 0 0 190 2
1385 1267
1297 1267
3 3 91 0 0 4224 0 74 73 0 0 4
1524 1472
1741 1472
1741 1392
1762 1392
3 2 92 0 0 4224 0 77 73 0 0 2
1521 1383
1763 1383
3 1 93 0 0 4224 0 80 73 0 0 4
1518 1282
1740 1282
1740 1374
1762 1374
0 3 85 0 0 0 0 0 75 190 0 3
1297 1464
1297 1512
1389 1512
0 3 85 0 0 4096 0 0 76 217 0 3
1297 1208
1297 1466
1388 1466
0 2 13 0 0 0 0 0 75 192 0 3
1282 1457
1282 1503
1389 1503
0 2 13 0 0 0 0 0 76 197 0 3
1282 1418
1282 1457
1388 1457
0 1 11 0 0 0 0 0 75 201 0 3
1217 1399
1217 1494
1389 1494
0 1 12 0 0 0 0 0 76 199 0 3
1254 1409
1254 1448
1388 1448
2 4 94 0 0 12416 0 74 75 0 0 4
1478 1481
1470 1481
1470 1503
1434 1503
4 1 95 0 0 4224 0 76 74 0 0 4
1433 1457
1469 1457
1469 1463
1478 1463
0 3 13 0 0 4096 0 0 78 215 0 3
1282 1200
1282 1418
1388 1418
0 3 88 0 0 0 0 0 79 208 0 3
1268 1316
1268 1368
1388 1368
0 2 12 0 0 0 0 0 78 207 0 3
1254 1307
1254 1409
1388 1409
0 2 83 0 0 0 0 0 79 222 0 3
1234 1097
1234 1359
1388 1359
0 1 11 0 0 0 0 0 78 202 0 3
1217 1346
1217 1400
1388 1400
0 1 11 0 0 0 0 0 79 220 0 3
1217 1142
1217 1350
1388 1350
4 2 96 0 0 4224 0 78 77 0 0 4
1433 1409
1466 1409
1466 1392
1475 1392
4 1 97 0 0 4224 0 79 77 0 0 4
1433 1359
1465 1359
1465 1374
1475 1374
4 2 98 0 0 4224 0 81 80 0 0 4
1432 1307
1457 1307
1457 1291
1472 1291
4 1 99 0 0 4224 0 82 80 0 0 4
1430 1258
1459 1258
1459 1273
1472 1273
0 2 12 0 0 4096 0 0 81 237 0 3
1254 932
1254 1307
1387 1307
0 3 88 0 0 0 0 0 81 209 0 3
1268 1256
1268 1316
1387 1316
0 2 88 0 0 0 0 0 82 219 0 3
1268 1156
1268 1258
1385 1258
0 1 84 0 0 0 0 0 81 211 0 3
1200 1249
1200 1298
1387 1298
0 1 84 0 0 0 0 0 82 216 0 3
1200 1189
1200 1249
1385 1249
4 3 100 0 0 4224 0 84 83 0 0 4
1428 1200
1758 1200
1758 1151
1767 1151
4 2 101 0 0 4224 0 85 83 0 0 4
1429 1153
1621 1153
1621 1142
1768 1142
3 1 102 0 0 4224 0 86 83 0 0 4
1429 1108
1757 1108
1757 1133
1767 1133
0 2 13 0 0 0 0 0 84 226 0 3
1282 1048
1282 1200
1383 1200
0 1 84 0 0 0 0 0 84 227 0 3
1200 1039
1200 1191
1383 1191
0 3 85 0 0 0 0 0 84 218 0 3
1297 1162
1297 1209
1383 1209
0 3 85 0 0 0 0 0 85 221 0 3
1297 1117
1297 1162
1384 1162
0 2 88 0 0 4096 0 0 85 239 0 4
1268 870
1268 1156
1384 1156
1384 1153
0 1 11 0 0 0 0 0 85 238 0 3
1217 921
1217 1144
1384 1144
0 2 85 0 0 0 0 0 86 225 0 3
1297 1057
1297 1117
1384 1117
0 1 83 0 0 0 0 0 86 229 0 3
1234 988
1234 1099
1384 1099
0 3 14 0 0 0 0 0 91 224 0 3
1316 890
1316 941
1383 941
0 3 14 0 0 4096 0 0 92 255 0 3
1316 619
1316 890
1381 890
0 3 85 0 0 4096 0 0 88 247 0 3
1297 785
1297 1057
1390 1057
0 2 13 0 0 0 0 0 88 228 0 3
1282 997
1282 1048
1390 1048
0 1 84 0 0 0 0 0 88 230 0 3
1200 979
1200 1039
1390 1039
0 3 13 0 0 4096 0 0 89 252 0 3
1282 717
1282 997
1388 997
0 2 83 0 0 0 0 0 89 248 0 3
1234 766
1234 988
1388 988
0 1 84 0 0 0 0 0 89 261 0 3
1200 547
1200 979
1388 979
3 3 103 0 0 4224 0 87 96 0 0 4
1512 1012
1751 1012
1751 914
1766 914
4 2 104 0 0 4224 0 88 87 0 0 3
1435 1048
1466 1048
1466 1021
4 1 105 0 0 4224 0 89 87 0 0 3
1433 988
1466 988
1466 1003
3 2 106 0 0 4224 0 90 96 0 0 3
1508 906
1767 906
1767 905
4 2 107 0 0 4224 0 91 90 0 0 3
1428 932
1462 932
1462 915
4 1 108 0 0 4224 0 92 90 0 0 3
1426 881
1462 881
1462 897
0 2 12 0 0 0 0 0 91 240 0 3
1254 881
1254 932
1383 932
0 1 11 0 0 0 0 0 91 246 0 3
1217 814
1217 923
1383 923
0 1 88 0 0 0 0 0 92 244 0 3
1268 832
1268 872
1381 872
0 2 12 0 0 0 0 0 92 245 0 3
1254 824
1254 881
1381 881
3 1 109 0 0 4224 0 93 96 0 0 4
1495 801
1750 801
1750 896
1766 896
3 1 110 0 0 4224 0 95 93 0 0 4
1419 776
1442 776
1442 792
1449 792
4 2 111 0 0 4224 0 94 93 0 0 4
1422 824
1443 824
1443 810
1449 810
0 3 88 0 0 4096 0 0 94 265 0 3
1268 469
1268 833
1377 833
0 2 12 0 0 0 0 0 94 254 0 3
1254 646
1254 824
1377 824
0 1 11 0 0 0 0 0 94 251 0 3
1217 702
1217 815
1377 815
0 2 85 0 0 0 0 0 95 264 0 3
1297 517
1297 785
1374 785
0 1 83 0 0 4224 0 0 95 270 0 3
1234 354
1234 767
1374 767
3 3 112 0 0 12416 0 99 97 0 0 4
1763 638
1723 638
1723 708
1553 708
3 2 113 0 0 4224 0 98 99 0 0 4
1552 655
1715 655
1715 629
1764 629
0 1 11 0 0 8192 0 0 97 266 0 4
1217 497
1217 702
1498 702
1498 699
2 0 13 0 0 0 0 97 0 0 253 3
1498 717
1282 717
1282 664
0 2 13 0 0 0 0 0 98 260 0 3
1282 557
1282 664
1497 664
0 1 12 0 0 0 0 0 98 299 0 3
1251 301
1251 646
1497 646
0 1 14 0 0 8320 0 0 99 259 0 3
1316 619
1316 620
1763 620
3 1 114 0 0 4224 0 104 106 0 0 4
1509 363
1734 363
1734 465
1768 465
3 2 115 0 0 4224 0 101 106 0 0 4
1503 494
1733 494
1733 474
1769 474
4 3 116 0 0 4224 0 100 106 0 0 4
1414 557
1763 557
1763 483
1768 483
0 3 14 0 0 0 0 0 100 298 0 5
1316 319
1316 619
1316 619
1316 566
1369 566
0 2 13 0 0 4096 0 0 100 296 0 3
1282 267
1282 557
1369 557
0 1 84 0 0 0 0 0 100 297 0 3
1200 259
1200 548
1369 548
3 2 117 0 0 4224 0 102 101 0 0 4
1415 508
1453 508
1453 503
1457 503
3 1 118 0 0 4224 0 103 101 0 0 3
1415 460
1457 460
1457 485
0 2 85 0 0 0 0 0 102 268 0 3
1297 462
1297 517
1370 517
0 2 88 0 0 0 0 0 103 269 0 3
1265 444
1265 469
1370 469
0 1 11 0 0 0 0 0 102 267 0 3
1217 497
1217 499
1370 499
0 1 11 0 0 0 0 0 103 301 0 5
1217 216
1217 497
1217 497
1217 451
1370 451
2 2 85 0 0 4224 0 124 105 0 0 5
1297 147
1297 462
1297 462
1297 417
1367 417
0 1 88 0 0 0 0 0 105 300 0 5
1265 234
1265 444
1265 444
1265 399
1367 399
1 2 83 0 0 0 0 104 122 0 0 3
1463 354
1234 354
1234 145
3 2 119 0 0 8320 0 105 104 0 0 3
1412 408
1412 372
1463 372
3 0 120 0 0 0 0 107 0 0 350 2
633 797
633 797
1 0 121 0 0 4096 0 108 0 0 282 2
242 1424
240 1424
4 0 122 0 0 4096 0 108 0 0 281 2
244 1459
244 1461
3 0 123 0 0 4096 0 108 0 0 277 2
244 1435
244 1438
2 0 124 0 0 0 0 108 0 0 278 2
244 1447
244 1447
0 0 123 0 0 8320 0 0 0 284 0 3
384 1298
384 1438
240 1438
0 0 124 0 0 8320 0 0 0 283 0 3
404 1386
404 1447
240 1447
0 4 122 0 0 4096 0 0 112 281 0 3
338 1461
338 1353
324 1353
0 1 121 0 0 4096 0 0 112 282 0 3
334 1209
334 1326
324 1326
3 0 122 0 0 4224 0 116 0 0 0 3
442 1461
240 1461
240 1456
3 0 121 0 0 8320 0 113 0 0 0 3
438 1209
240 1209
240 1429
3 3 124 0 0 0 0 115 112 0 0 4
441 1386
366 1386
366 1344
324 1344
3 2 123 0 0 0 0 114 112 0 0 4
439 1298
369 1298
369 1335
324 1335
2 13 125 0 0 8320 0 116 131 0 0 4
497 1470
1117 1470
1117 466
1080 466
2 12 126 0 0 8320 0 115 131 0 0 4
496 1395
1128 1395
1128 457
1080 457
2 11 127 0 0 8320 0 114 131 0 0 4
494 1307
1136 1307
1136 448
1080 448
2 10 128 0 0 8320 0 113 131 0 0 4
493 1218
1144 1218
1144 439
1080 439
1 1 129 0 0 4224 0 117 116 0 0 3
687 1107
687 1452
497 1452
2 1 130 0 0 4224 0 117 115 0 0 3
681 1107
681 1377
496 1377
3 1 131 0 0 4224 0 117 114 0 0 3
675 1107
675 1289
494 1289
4 1 132 0 0 8320 0 117 113 0 0 3
669 1107
669 1200
493 1200
1 0 18 0 0 0 0 135 0 0 294 3
803 597
803 713
900 713
1 6 18 0 0 0 0 127 137 0 0 4
907 528
900 528
900 783
840 783
0 3 14 0 0 0 0 0 119 298 0 3
1316 280
1638 280
1638 277
0 2 13 0 0 12416 0 0 119 307 0 4
1265 33
1282 33
1282 268
1638 268
2 1 84 0 0 0 0 125 119 0 0 3
1200 145
1200 259
1638 259
0 2 14 0 0 0 0 0 120 308 0 4
1297 22
1316 22
1316 319
1636 319
0 1 12 0 0 12288 0 0 120 306 0 4
1234 42
1251 42
1251 301
1636 301
2 2 88 0 0 8320 0 123 118 0 0 3
1265 147
1265 234
1638 234
0 1 11 0 0 12288 0 0 118 305 0 4
1198 54
1217 54
1217 216
1638 216
3 3 133 0 0 4224 0 120 121 0 0 3
1691 310
1765 310
1765 272
4 2 134 0 0 4224 0 119 121 0 0 3
1683 268
1766 268
1766 263
3 1 135 0 0 4224 0 118 121 0 0 3
1683 225
1765 225
1765 254
0 1 11 0 0 0 0 0 125 321 0 6
1009 299
1009 232
1041 232
1041 54
1200 54
1200 109
1 0 12 0 0 0 0 122 0 0 320 5
1234 109
1234 40
1032 40
1032 222
996 222
1 0 13 0 0 0 0 123 0 0 319 5
1265 111
1265 32
1024 32
1024 212
985 212
0 1 14 0 0 0 0 0 124 318 0 5
972 201
1014 201
1014 22
1297 22
1297 111
1 0 12 0 0 0 0 142 0 0 320 2
835 112
835 182
1 9 136 0 0 8320 0 1 131 0 0 3
1007 499
1007 493
1016 493
1 0 15 0 0 0 0 130 0 0 340 3
906 423
860 423
860 651
1 0 16 0 0 0 0 128 0 0 339 3
906 457
870 457
870 660
1 0 17 0 0 0 0 129 0 0 338 3
906 490
880 490
880 669
2 8 137 0 0 8320 0 127 131 0 0 4
943 528
969 528
969 475
1016 475
2 7 138 0 0 12416 0 129 131 0 0 4
942 490
962 490
962 466
1016 466
2 6 139 0 0 4224 0 128 131 0 0 2
942 457
1016 457
2 5 140 0 0 12416 0 130 131 0 0 4
942 423
957 423
957 448
1016 448
0 4 14 0 0 0 0 0 131 356 0 4
941 161
972 161
972 439
1016 439
0 3 13 0 0 0 0 0 131 355 0 5
882 172
882 174
985 174
985 430
1016 430
0 2 12 0 0 4224 0 0 131 367 0 6
400 182
835 182
835 184
996 184
996 421
1016 421
0 1 11 0 0 0 0 0 131 354 0 4
867 299
1009 299
1009 412
1016 412
0 0 141 0 0 4096 0 0 0 330 347 3
78 205
78 821
252 821
5 0 141 0 0 0 0 149 0 0 330 2
617 204
617 205
1 0 142 0 0 0 0 149 0 0 329 2
617 279
617 279
5 0 141 0 0 0 0 148 0 0 330 2
441 204
441 205
1 0 142 0 0 4096 0 148 0 0 329 4
441 279
441 278
441 278
441 279
5 0 141 0 0 0 0 147 0 0 330 2
253 204
253 205
1 0 142 0 0 0 0 147 0 0 329 2
253 279
253 279
1 1 142 0 0 8320 0 153 2 0 0 5
788 280
788 279
253 279
253 281
166 281
5 0 141 0 0 4224 0 153 0 0 0 2
788 205
75 205
0 3 17 0 0 0 0 0 137 332 0 3
774 784
774 801
792 801
1 0 17 0 0 0 0 137 0 0 338 3
792 783
792 784
774 784
1 0 15 0 0 0 0 139 0 0 334 2
469 770
435 770
3 0 15 0 0 0 0 139 0 0 340 3
469 788
435 788
435 761
1 0 17 0 0 0 0 134 0 0 338 2
775 597
775 669
1 0 16 0 0 0 0 133 0 0 339 2
730 596
730 660
1 0 15 0 0 0 0 132 0 0 340 2
687 597
687 651
6 0 17 0 0 0 0 138 0 0 0 4
730 784
774 784
774 669
897 669
6 0 16 0 0 0 0 139 0 0 0 4
517 770
664 770
664 660
897 660
6 0 15 0 0 0 0 140 0 0 0 4
405 761
435 761
435 651
897 651
2 0 2 0 0 0 0 138 0 0 343 3
675 793
664 793
664 866
2 0 2 0 0 0 0 139 0 0 343 3
462 779
458 779
458 866
2 2 2 0 0 12288 0 140 137 0 0 6
350 770
322 770
322 866
770 866
770 792
785 792
4 0 141 0 0 0 0 138 0 0 347 3
706 832
706 837
700 837
4 0 141 0 0 0 0 139 0 0 347 2
493 818
493 837
4 0 141 0 0 0 0 140 0 0 347 4
381 809
381 829
357 829
357 837
1 4 141 0 0 0 0 136 137 0 0 4
252 764
252 837
816 837
816 831
1 3 141 0 0 0 0 136 140 0 0 3
252 764
252 779
357 779
1 1 141 0 0 0 0 136 140 0 0 3
252 764
252 761
357 761
0 3 120 0 0 12416 0 0 138 0 0 4
629 797
655 797
655 802
682 802
0 1 143 0 0 4224 0 0 138 0 0 4
629 797
660 797
660 784
682 784
5 2 144 0 0 16512 0 140 107 0 0 7
411 779
411 797
458 797
458 823
569 823
569 806
584 806
5 1 145 0 0 4224 0 139 107 0 0 2
523 788
584 788
1 7 11 0 0 20608 0 141 147 0 0 8
790 106
819 106
819 214
867 214
867 299
209 299
209 252
229 252
1 0 13 0 0 0 0 143 0 0 370 5
883 113
883 166
882 166
882 174
639 174
1 0 14 0 0 0 0 144 0 0 371 6
935 113
941 113
941 161
930 161
930 136
726 136
3 0 2 0 0 0 0 147 0 0 360 4
283 243
283 313
284 313
284 328
3 0 2 0 0 0 0 148 0 0 360 2
471 243
471 328
3 0 2 0 0 0 0 149 0 0 360 2
647 243
647 328
0 3 2 0 0 41088 0 0 153 343 0 13
531 866
531 914
173 914
173 542
480 542
480 425
426 425
426 349
208 349
208 328
825 328
825 244
818 244
1 2 146 0 0 12416 0 3 145 0 0 4
172 498
196 498
196 436
287 436
3 1 147 0 0 8336 0 146 145 0 0 4
154 390
154 381
287 381
287 418
4 0 148 0 0 8320 0 151 0 0 364 3
298 104
293 104
293 253
4 2 148 0 0 0 0 147 147 0 0 6
277 234
323 234
323 253
293 253
293 252
277 252
3 0 14 0 0 0 0 151 0 0 371 3
343 95
657 95
657 135
0 2 13 0 0 0 0 0 151 370 0 4
642 165
419 165
419 104
343 104
7 1 12 0 0 0 0 148 151 0 0 4
417 252
400 252
400 113
343 113
3 0 149 0 0 8320 0 152 0 0 369 3
568 144
487 144
487 249
4 2 149 0 0 0 0 148 148 0 0 6
465 234
515 234
515 249
487 249
487 252
465 252
7 1 13 0 0 0 0 149 152 0 0 6
593 252
574 252
574 174
642 174
642 153
613 153
0 2 14 0 0 0 0 0 152 373 0 3
726 235
726 135
613 135
2 0 14 0 0 0 0 149 0 0 373 4
641 252
711 252
711 253
726 253
4 7 14 0 0 0 0 149 153 0 0 4
641 234
726 234
726 253
764 253
0 1 150 0 0 4096 0 0 150 375 0 3
871 244
925 244
925 235
4 2 150 0 0 4224 0 153 153 0 0 4
812 235
871 235
871 253
812 253
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1030 658 1115 682
1040 666 1104 682
8 overflow
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
427 1558 528 1582
437 1566 517 1582
10 OPERANDO 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
176 1554 277 1578
186 1562 266 1578
10 OPERANDO 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1028 346 1073 370
1038 354 1062 370
3 ULA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
117 75 194 99
127 83 183 99
7 PASSO 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
117 57 282 81
127 65 271 81
18 CONTADOR CRESCENTE
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
581 613 634 637
591 621 623 637
4 LFSR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
276 1162 377 1186
286 1170 366 1186
10 COMPARADOR
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
602 1006 743 1030
612 1014 732 1030
15 ENTRADA USU�RIO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
328 1616 373 1640
338 1624 362 1640
3 ___
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
